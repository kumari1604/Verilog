`timescale 1ns / 1ps



module decoder_enable(
    input en,
    input [1:0] x,
    output [3:0] y
    );
    wire x1_bar,x0_bar;               // if enable=0 y0=y1=y2=y3=0
	                                   // if enable=1 y0=x1'x0', y1=x1'x0 , y2=x1x0' , y3=x1x0
    not(x1_bar,x[1]);
    not(x0_bar,x[0]);
    and(y[0],x1_bar,x0_bar,en);
    and(y[1],x1_bar,x[0],en);
    and(y[2],x[1],x0_bar,en);
    and(y[3],x[1],x[0],en);
endmodule
